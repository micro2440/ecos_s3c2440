# ====================================================================
#
#      gfx_png.cdl
#
#      libpng configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Alexander Neundorf <neundorf@kde.org>
# Contributors:
# Date:           2008-03-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_GFX_PNG {
    display       "PNG library"
    description   "
                  This package provides support for compression and
                  decompression."
#    include_dir   cyg/png 

    requires      CYGPKG_ISOINFRA
    requires      CYGPKG_COMPRESS_ZLIB
    requires      CYGPKG_CRC
    requires      CYGPKG_LIBC_SETJMP

    compile       png.c pngset.c pngget.c pngrutil.c pngtrans.c pngwutil.c 
    compile       pngread.c pngrio.c pngwio.c pngwrite.c pngrtran.c 
    compile       pngwtran.c pngmem.c pngerror.c pngread.c

#    cdl_interface CYGINT_COMPRESS_ZLIB_LOCAL_ALLOC {
#        display "Override memory allocation routines."
#    }

     cdl_option CYGFUN_PNG_WITH_STDIO {
        display "With file (stdio) functions"
        default_value 0
        requires CYGPKG_IO_FILEIO
     }

     cdl_option CYGFUN_PNG_NO_WRITE {
        display "Disable writing function"
        default_value 0
     }

     cdl_option CYGFUN_PNG_NO_READ {
        display "Disable reading function"
        default_value 0
     }


    cdl_component CYGPKG_GFX_PNG_OPTIONS {
        display "PNG compress and decompress package build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."

        cdl_option CYGPKG_GFX_PNG_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D__ECOS__ -O3 -funroll-loops" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in addition
                to the set of global flags."
        }
    }
 

}

# ====================================================================
# EOF compress_zlib.cdl
