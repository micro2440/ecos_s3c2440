# ====================================================================
#
#      pwin.cdl
#
#      eCos PW graphic library configuration data 
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2004 Savin Zlobec
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s): Savin Zlobec 
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_PWIN {
    display       "PW graphic library" 
    description   "PW graphic library."
    
    compile             \
        pw_display.c    \
        pw_init.c       \
        pw_window.c     \
        pw_region.c     \
        pw_rgalloc.c    \
        pw_draw.c       \
        pw_bitmap.c     \
        pw_event.c      \
        pw_timeout.c    \
        pw_diag.c

    cdl_option CYGBLD_PWIN_SYNTH_DRIVER {
        display       "PW graphic library synth target display driver"
        active_if     CYGPKG_HAL_SYNTH
        default_value 1
        compile       drivers/dd_synth.c    
    }

    cdl_component CYGPKG_PWIN_OPTIONS {
        display "PW graphic library build options"
        flavor  none
        description   "
	        Package specific build options including control over
	        compiler flags used only in building this package,
	        and details of which tests are built."

        cdl_option CYGPKG_PWIN_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in 
                addition to the set of global flags."
        }

        cdl_option CYGPKG_PWIN_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_PWIN_TESTS {
            display     "PW graphic library tests"
            flavor      data
            no_define
            calculated  { "tests/pw_test" }
            description "
                This option specifies the set of tests for the PW 
                graphic library."
        }
    }
}

# EOF pwin.cdl
